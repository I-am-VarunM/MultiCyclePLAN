module SBOX(bb_in7, bb_in6, bb_in5, bb_in4, bb_in3, bb_in2, bb_in1, bb_in0, bb_out7, bb_out6, bb_out5, bb_out4, bb_out3, bb_out2, bb_out1, bb_out0);
  input bb_in7, bb_in6, bb_in5, bb_in4, bb_in3, bb_in2, bb_in1, bb_in0;
  output bb_out7, bb_out6, bb_out5, bb_out4, bb_out3, bb_out2, bb_out1, bb_out0;
  wire bb_in7, bb_in6, bb_in5, bb_in4, bb_in3, bb_in2, bb_in1, bb_in0;
  wire bb_out7, bb_out6, bb_out5, bb_out4, bb_out3, bb_out2, bb_out1, bb_out0;
  wire n_7, n_9, n_20, n_24, n_25, n_26, n_30, n_31;
  wire n_36, n_43, n_45, n_46, n_51, n_52, n_53, n_54;
  wire n_55, n_56, n_58, n_59, n_65, n_69, n_71, n_77;
  wire n_84, n_86, n_87, n_91, n_92, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_103, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_117, n_119, n_123;
  wire n_124, n_126, n_127, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_141, n_142, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_153, n_155;
  wire n_156, n_163, n_164, n_168, n_169, n_174, n_176, n_178;
  wire n_181, n_182, n_183, n_184, n_185, n_189, n_192, n_193;
  wire n_194, n_196, n_198, n_199, n_200, n_201, n_204, n_205;
  wire n_206, n_207, n_208, n_209, n_212, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_229, n_230, n_231, n_232, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_245;
  wire n_246, n_248, n_249, n_250, n_251, n_252, n_253, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_264, n_265, n_266;
  wire n_267, n_269, n_270, n_274, n_275, n_276, n_277, n_279;
  wire n_280, n_281, n_282, n_283, n_284, n_286, n_287, n_291;
  wire n_292, n_293, n_294, n_296, n_298, n_299, n_300, n_301;
  wire n_302, n_303, n_304, n_306, n_307, n_308, n_309, n_311;
  wire n_312, n_314, n_334, n_335, n_336, n_337, n_338, n_342;
  wire n_343, n_346, n_408, n_409, n_412, n_413, n_414, n_416;
  wire n_417, n_418, n_419, n_429, n_430, n_461, n_462, n_463;
  wire n_464, n_465, n_466, n_472, n_473, n_474, n_475, n_476;
  wire n_478, n_479, n_480, n_481, n_518, n_519, n_521, n_522;
  wire n_523, n_544, n_545, n_547, n_548, n_549, n_550, n_552;
  wire n_553, n_554, n_559, n_560, n_561, n_562, n_563, n_565;
  wire n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573;
  wire n_574, n_575, n_578, n_579, n_580, n_581, n_582, n_583;
  wire n_584, n_585, n_586, n_587, n_588, n_589, n_590, n_591;
  wire n_607, n_609, n_612, n_613, n_614, n_615, n_647, n_648;
  wire n_649, n_650, n_651, n_652, n_654, n_655;
  xnor XNOR2_182 (n_25, bb_in0, bb_in1);
  not NOT1_183 (n_9, bb_in1);
  xor XOR2_186 (n_336, bb_in1, bb_in2);
  xnor XNOR2_194 (n_412, bb_in6, bb_in7);
  not NOT1_197 (n_413, bb_in6);
  not NOT1_199 (n_7, bb_in7);
  xor XOR2_214 (n_475, bb_in6, bb_in4);
  not NOT1_218 (n_479, bb_in4);
  xor XOR2_225 (n_544, bb_in4, bb_in2);
  not NOT1_228 (n_547, bb_in2);
  not NOT1_230 (n_549, bb_in3);
  xor XOR2_231 (n_553, bb_in1, bb_in5);
  not NOT1_232 (n_554, bb_in5);
  not NOT1_179 (n_26, n_25);
  nand NAND2_196 (n_414, n_413, bb_in7);
  nand NAND2_216 (n_478, n_413, bb_in4);
  nand NAND2_180 (n_24, n_7, bb_in5);
  nand NAND2_198 (n_416, n_7, bb_in6);
  xnor XNOR2_213 (n_476, n_475, n_553);
  nand NAND2_217 (n_480, n_479, bb_in6);
  xnor XNOR2_224 (n_545, n_544, bb_in3);
  nand NAND2_227 (n_548, n_547, bb_in3);
  nand NAND2_229 (n_550, n_549, bb_in2);
  nand NAND2_181 (n_20, n_554, bb_in7);
  nand NAND2_195 (n_417, n_414, n_416);
  nand NAND2_215 (n_481, n_478, n_480);
  nand NAND2_178 (n_30, n_24, n_20);
  not NOT1_173 (n_45, n_476);
  nand NAND2_211 (n_472, n_548, n_550);
  nand NAND2_270 (n_647, n_548, n_550);
  nand NAND2_168 (n_55, n_545, n_417);
  xnor XNOR2_265 (n_607, n_336, n_417);
  xnor XNOR2_175 (n_98, n_9, n_481);
  not NOT1_177 (n_31, n_30);
  xnor XNOR2_212 (n_474, n_472, n_30);
  not NOT1_170 (n_54, n_45);
  xnor XNOR2_226 (n_552, n_479, n_647);
  xnor XNOR2_272 (n_648, bb_in7, n_647);
  xnor XNOR2_275 (n_651, bb_in7, n_647);
  nor NOR2_219 (n_518, n_607, n_476);
  not NOT1_264 (n_84, n_607);
  not NOT1_203 (n_430, n_98);
  not NOT1_176 (n_36, n_31);
  not NOT1_172 (n_52, n_474);
  not NOT1_158 (n_65, n_54);
  xnor XNOR2_210 (n_473, n_472, n_54);
  nand NAND2_169 (n_46, n_552, n_412);
  not NOT1_271 (n_649, n_648);
  xnor XNOR2_273 (n_650, bb_in6, n_648);
  nand NAND2_274 (n_652, n_651, n_26);
  not NOT1_263 (n_609, n_84);
  nand NAND2_268 (n_614, n_84, n_36);
  xnor XNOR2_269 (n_615, n_98, n_84);
  nor NOR2_163 (n_71, n_430, n_54);
  nor NOR2_166 (n_58, n_474, n_430);
  nor NOR2_167 (n_56, n_31, n_430);
  not NOT1_202 (n_429, n_430);
  not NOT1_174 (n_43, n_36);
  nand NAND2_220 (n_519, n_650, n_36);
  not NOT1_162 (n_53, n_52);
  not NOT1_156 (n_100, n_65);
  nand NAND2_161 (n_204, n_55, n_46);
  nand NAND2_165 (n_59, n_649, n_25);
  nand NAND2_159 (n_77, n_650, n_45);
  not NOT1_188 (n_337, n_650);
  nor NOR2_164 (n_69, n_53, n_609);
  xnor XNOR2_150 (n_95, n_58, n_615);
  xnor XNOR2_143 (n_106, n_56, n_77);
  xnor XNOR2_146 (n_201, n_53, n_429);
  nand NAND2_147 (n_99, n_204, n_429);
  nand NAND2_145 (n_103, n_84, n_43);
  not NOT1_171 (n_51, n_43);
  xnor XNOR2_193 (n_408, n_518, n_519);
  xnor XNOR2_223 (n_521, n_31, n_519);
  nor NOR2_155 (n_86, n_53, n_337);
  nand NAND2_152 (n_92, n_204, n_54);
  not NOT1_157 (n_221, n_204);
  nand NAND2_266 (n_612, n_204, n_84);
  nand NAND2_160 (n_110, n_652, n_59);
  nand NAND2_134 (n_119, n_337, n_65);
  not NOT1_187 (n_338, n_337);
  xnor XNOR2_127 (n_139, n_69, n_106);
  xnor XNOR2_192 (n_409, n_95, n_408);
  not NOT1_138 (n_229, n_201);
  nand NAND2_153 (n_91, n_609, n_51);
  xnor XNOR2_222 (n_522, n_518, n_521);
  nand NAND2_139 (n_111, n_110, n_221);
  nor NOR2_141 (n_108, n_221, n_337);
  nand NAND2_142 (n_107, n_221, n_65);
  xnor XNOR2_267 (n_613, n_84, n_221);
  xnor XNOR2_133 (n_123, n_614, n_612);
  xnor XNOR2_137 (n_112, n_110, n_473);
  nand NAND2_144 (n_105, n_110, n_204);
  nand NAND2_148 (n_97, n_110, n_52);
  nand NAND2_149 (n_96, n_110, n_36);
  nand NAND2_151 (n_94, n_110, n_65);
  not NOT1_154 (n_87, n_110);
  nand NAND2_136 (n_117, n_338, n_54);
  xnor XNOR2_115 (n_149, n_99, n_139);
  nand NAND2_135 (n_217, n_91, n_103);
  xnor XNOR2_125 (n_131, n_94, n_108);
  nand NAND2_129 (n_134, n_92, n_107);
  xnor XNOR2_123 (n_135, n_86, n_613);
  xnor XNOR2_128 (n_127, n_337, n_105);
  xnor XNOR2_131 (n_126, n_337, n_97);
  xnor XNOR2_132 (n_124, n_71, n_96);
  nand NAND2_140 (n_109, n_87, n_204);
  nand NAND2_126 (n_227, n_119, n_117);
  not NOT1_109 (n_150, n_149);
  xnor XNOR2_118 (n_145, n_131, n_409);
  xnor XNOR2_120 (n_156, n_112, n_134);
  xor XOR2_277 (n_654, n_614, n_134);
  not NOT1_119 (n_136, n_135);
  xnor XNOR2_116 (n_147, n_127, n_139);
  xnor XNOR2_221 (n_523, n_126, n_522);
  xnor XNOR2_121 (n_137, n_123, n_124);
  nand NAND2_130 (n_207, n_109, n_111);
  not NOT1_122 (n_133, n_227);
  not NOT1_111 (n_146, n_145);
  nand NAND2_246 (n_571, n_145, n_654);
  xnor XNOR2_105 (n_174, n_156, n_147);
  not NOT1_114 (n_141, n_654);
  not NOT1_110 (n_148, n_147);
  nand NAND2_107 (n_153, n_523, n_149);
  not NOT1_112 (n_144, n_523);
  nand NAND2_113 (n_142, n_137, n_135);
  not NOT1_117 (n_138, n_137);
  not NOT1_124 (n_132, n_207);
  nand NAND2_245 (n_570, n_146, n_141);
  xnor XNOR2_103 (n_164, n_156, n_148);
  nand NAND2_106 (n_155, n_144, n_150);
  nand NAND2_108 (n_151, n_138, n_136);
  nand NAND2_244 (n_572, n_570, n_571);
  nand NAND2_255 (n_584, n_155, n_153);
  nand NAND2_104 (n_163, n_151, n_142);
  not NOT1_243 (n_573, n_572);
  nand NAND3_248 (n_575, n_572, n_584, n_164);
  nand NAND2_253 (n_582, n_572, n_163);
  nand NAND2_101 (n_178, n_584, n_174);
  not NOT1_257 (n_585, n_584);
  not NOT1_260 (n_588, n_584);
  not NOT1_102 (n_168, n_163);
  nand NAND3_98 (n_169, n_584, n_573, n_168);
  nand NAND2_99 (n_183, n_573, n_163);
  not NOT1_251 (n_579, n_573);
  not NOT1_201 (n_419, n_575);
  nor NOR2_97 (n_181, n_178, n_582);
  not NOT1_191 (n_346, n_178);
  nand NAND2_237 (n_561, n_178, n_168);
  nand NAND4_256 (n_586, n_585, n_572, n_174, n_163);
  nand NAND3_258 (n_587, n_585, n_572, n_168);
  nand NAND3_261 (n_590, n_588, n_164, n_163);
  nand NAND2_262 (n_591, n_588, n_164);
  nand NAND3_100 (n_176, n_584, n_174, n_168);
  nor NOR2_247 (n_574, n_572, n_168);
  nand NAND3_249 (n_578, n_168, n_174, n_572);
  nand NAND2_252 (n_581, n_572, n_168);
  nand NAND2_92 (n_192, n_591, n_169);
  nor NOR2_93 (n_189, n_174, n_183);
  nand NAND2_95 (n_184, n_183, n_581);
  nor NOR2_250 (n_580, n_579, n_591);
  nor NOR2_254 (n_583, n_178, n_579);
  nand NAND2_236 (n_560, n_346, n_574);
  nand NAND2_91 (n_193, n_586, n_176);
  not NOT1_96 (n_182, n_587);
  nand NAND2_94 (n_185, n_590, n_578);
  nand NAND2_259 (n_589, n_574, n_588);
  nor NOR2_88 (n_198, n_192, n_182);
  nor NOR2_89 (n_196, n_181, n_189);
  nand NAND2_90 (n_194, n_184, n_164);
  nor NOR2_235 (n_559, n_419, n_580);
  nor NOR2_87 (n_199, n_583, n_193);
  nand NAND3_200 (n_418, n_575, n_176, n_589);
  nand NAND2_84 (n_225, n_198, n_196);
  nand NAND2_85 (n_214, n_199, n_194);
  nand NAND3_234 (n_562, n_559, n_560, n_561);
  nor NOR2_86 (n_220, n_185, n_418);
  nand NAND2_67 (n_226, n_225, n_52);
  nand NAND2_68 (n_224, n_225, n_65);
  nand NAND2_69 (n_223, n_225, n_207);
  nand NAND2_73 (n_251, n_225, n_217);
  nand NAND2_74 (n_253, n_225, n_51);
  not NOT1_82 (n_200, n_225);
  nand NAND2_185 (n_334, n_225, n_204);
  nand NAND2_207 (n_462, n_225, n_227);
  nand NAND2_75 (n_216, n_214, n_227);
  nand NAND2_76 (n_215, n_214, n_201);
  nand NAND2_77 (n_212, n_214, n_36);
  nand NAND2_78 (n_209, n_214, n_52);
  nand NAND2_79 (n_208, n_214, n_207);
  nand NAND2_80 (n_206, n_214, n_65);
  nand NAND2_81 (n_205, n_214, n_204);
  nand NAND2_206 (n_461, n_214, n_217);
  not NOT1_233 (n_563, n_562);
  nand NAND2_238 (n_565, n_562, n_201);
  nor NOR2_66 (n_230, n_229, n_220);
  nor NOR2_70 (n_222, n_221, n_220);
  nor NOR2_71 (n_219, n_53, n_220);
  nor NOR2_72 (n_218, n_132, n_220);
  not NOT1_83 (n_238, n_220);
  xnor XNOR2_51 (n_276, n_212, n_224);
  xnor XNOR2_50 (n_252, n_223, n_251);
  xor XOR2_184 (n_335, n_334, n_253);
  nor NOR2_56 (n_241, n_229, n_200);
  xnor XNOR2_205 (n_463, n_461, n_462);
  xnor XNOR2_209 (n_465, n_461, n_462);
  xnor XNOR2_53 (n_249, n_208, n_230);
  xnor XNOR2_54 (n_248, n_205, n_219);
  nor NOR2_59 (n_237, n_133, n_563);
  nor NOR2_63 (n_232, n_43, n_563);
  nor NOR2_64 (n_231, n_100, n_563);
  not NOT1_240 (n_566, n_563);
  xnor XNOR2_52 (n_250, n_565, n_218);
  nand NAND2_57 (n_240, n_238, n_65);
  nand NAND2_58 (n_239, n_238, n_227);
  nand NAND2_60 (n_236, n_238, n_36);
  nand NAND2_61 (n_235, n_238, n_217);
  xnor XNOR2_38 (n_267, n_232, n_335);
  xnor XNOR2_208 (n_466, n_250, n_465);
  xnor XNOR2_47 (n_258, n_251, n_237);
  xnor XNOR2_48 (n_257, n_253, n_231);
  nand NAND2_239 (n_567, n_566, n_207);
  not NOT1_241 (n_568, n_566);
  nand NAND2_242 (n_569, n_566, n_217);
  xnor XNOR2_45 (n_260, n_209, n_240);
  xnor XNOR2_44 (n_261, n_215, n_239);
  xnor XNOR2_49 (n_256, n_206, n_236);
  xnor XNOR2_46 (n_259, n_216, n_235);
  xnor XNOR2_27 (n_306, n_260, n_267);
  xnor XNOR2_35 (n_280, n_567, n_466);
  xnor XNOR2_41 (n_266, n_249, n_258);
  xnor XNOR2_42 (n_265, n_248, n_257);
  not NOT1_55 (n_245, n_567);
  nor NOR2_62 (n_234, n_53, n_568);
  nor NOR2_65 (n_246, n_221, n_568);
  xnor XNOR2_43 (n_264, n_569, n_252);
  xnor XNOR2_40 (n_270, n_226, n_256);
  xnor XNOR2_39 (n_274, n_241, n_259);
  not NOT1_23 (n_312, n_306);
  not NOT1_29 (n_281, n_280);
  xnor XNOR2_204 (n_464, n_463, n_266);
  xnor XNOR2_33 (n_283, n_276, n_265);
  xnor XNOR2_278 (n_655, n_270, n_246);
  xnor XNOR2_36 (n_296, n_261, n_264);
  xnor XNOR2_32 (n_277, n_222, n_270);
  xnor XNOR2_31 (n_286, n_466, n_274);
  nand NAND2_34 (n_275, n_274, n_567);
  not NOT1_37 (n_269, n_274);
  xnor XNOR2_19 (n_293, n_464, n_280);
  not NOT1_190 (n_343, n_464);
  xnor XNOR2_21 (n_291, n_234, n_283);
  not NOT1_26 (n_284, n_283);
  nand NAND2_17 (n_298, n_655, n_296);
  not NOT1_22 (n_302, n_655);
  xnor XNOR2_16 (n_299, n_296, n_306);
  not NOT1_28 (n_282, n_296);
  xor XOR2_20 (n_292, n_276, n_277);
  not NOT1_25 (n_287, n_286);
  nand NAND2_30 (n_279, n_269, n_245);
  xnor XNOR2_8 (n_309, n_306, n_293);
  nand NAND2_18 (n_294, n_286, n_343);
  not NOT1_189 (n_342, n_343);
  xnor XNOR2_9 (n_308, n_291, n_292);
  xnor XNOR2_14 (n_301, n_284, n_655);
  nand NAND2_13 (n_303, n_302, n_282);
  xor XOR2_276 (bb_out6, n_302, n_312);
  nand NAND2_24 (bb_out3, n_279, n_275);
  xnor XNOR2_2 (bb_out4, n_301, n_309);
  xnor XNOR2_12 (n_304, n_342, bb_out3);
  nand NAND2_15 (n_300, n_287, n_342);
  nand NAND2_7 (n_311, n_303, n_298);
  xnor XNOR2_11 (n_307, n_306, bb_out3);
  xnor XNOR2_6 (bb_out1, n_312, n_304);
  nand NAND2_10 (n_314, n_300, n_294);
  xnor XNOR2_1 (bb_out2, n_281, n_311);
  xnor XNOR2_3 (bb_out0, n_307, n_308);
  xnor XNOR2_4 (bb_out7, n_299, n_314);
  xnor XNOR2_5 (bb_out5, n_312, n_314);

endmodule

module  Oracle (a, k, enca);
  input [7:0] a;
  input [7:0] k;
  output [7:0] enca;
  assign enca[7:0] = a[7:0] ^ k[7:0];
endmodule

module top;
reg [7:0]a;
reg [7:0] k;
wire [7:0] enca;
wire [7:0] out;
Oracle o1 (.a(a), .k(k), .enca(enca));
SBOX s1(.bb_in7(a[7]), .bb_in6(a[6]), .bb_in5(a[5]), .bb_in4(a[4]), .bb_in3(a[3]), .bb_in2(a[2]), .bb_in1(a[1]), .bb_in0(a[0]), .bb_out7(out[7]), .bb_out6(out[6]), .bb_out5(out[5]), .bb_out4(out[4]), .bb_out3(out[3]), .bb_out2(out[2]), .bb_out1(out[1]), .bb_out0(out[0]));
initial begin 
  a= 1;
  k = 8'b 10000000;
  $dumpfile(" 1.vcd");
	$dumpvars;
end
endmodule